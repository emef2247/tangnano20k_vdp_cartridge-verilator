// -----------------------------------------------------------------------------
//	tangnano20k_vdp_cartridge.v
//	Copyright (C)2025 Takayuki Hara (HRA!)
//	Modified 2026-01-02 by @emef2247 (Verilator integration)
//	Updated: restored proper rdata_en wiring and added guarded debug monitors
// -----------------------------------------------------------------------------

module tangnano20k_vdp_cartridge (
	input			clk,			//	PIN04		(27MHz)
	input			clk14m,			//	PIN80
	input			slot_reset_n,	//	PIN86
	input			slot_iorq_n,	//	PIN18
	input			slot_rd_n,		//	PIN15
	input			slot_wr_n,		//	PIN16
	output			slot_wait,		//	PIN72
	output			slot_intr,		//	PIN71
	output			slot_data_dir,	//	PIN19
	input	[7:0]	slot_a,			//	PIN17, 49, 48, 41, 42, 76, 31, 30
	inout	[7:0]	slot_d,			//	PIN73, 74, 75, 85, 77, 27, 28, 29
	output			oe_n,			//	PIN20
	input	[1:0]	dipsw,			//	PIN52, 53
	output			ws2812_led,		//	PIN79
	input	[1:0]	button,			//	PIN87, 88	KEY2, KEY1

	//	HDMI
	output			tmds_clk_p,		//	(PIN33/34)
	output			tmds_clk_n,		//	dummy
	output	[2:0]	tmds_d_p,		//	(PIN39/40), (PIN37/38), (PIN35/36)
	output	[2:0]	tmds_d_n,		//	dummy

	output			O_sdram_clk,
	output			O_sdram_cke,
	output			O_sdram_cs_n,	// chip select
	output			O_sdram_ras_n,	// row address select
	output			O_sdram_cas_n,	// columns address select
	output			O_sdram_wen_n,	// write enable
	inout	[31:0]	IO_sdram_dq,	// 32 bit bidirectional data bus
	output	[10:0]	O_sdram_addr,	// 11 bit multiplexed address bus
	output	[ 1:0]	O_sdram_ba,		// two banks
	output	[ 3:0]	O_sdram_dqm,	// data mask

	// --------------------------------------------------------------------
	// [MOD] Raw video output from VDP core (for Verilator / openMSX)
	// --------------------------------------------------------------------
    output          display_hs,
    output          display_vs,
    output          display_en,
    output  [7:0]   display_r,
    output  [7:0]   display_g,
    output  [7:0]   display_b,
	
	// --------------------------------------------------------------------
	// [MOD] Debug/functional VRAM bus exported from VDP core.
	// --------------------------------------------------------------------
	output	[17:0]	dbg_vram_address,
	output	[31:0]	dbg_vram_wdata,
	input	[31:0]	dbg_vram_rdata,
	output			dbg_vram_valid,
	output			dbg_vram_write,
	output			dbg_vram_rdata_en
);
	reg				ff_reset_n0 = 1'b0;
	reg				ff_reset_n1 = 1'b0;
	reg				ff_reset_n2_1 = 1'b0;
	reg				ff_reset_n2_2 = 1'b0;
	wire			pll_lock215;
	wire			pll_lock85;
	wire			clk42m;				//	42.95454MHz
	wire			clk85m;				//	85.90908MHz
	wire			clk85m_n;			//	85.90908MHz (180deg phase shift)
	wire			clk215m;			//	214.7727MHz
	wire			reset_n;
	wire			reset_n2;
	wire	[2:0]	w_bus_address;
	wire			w_bus_ioreq;
	wire			w_bus_write;
	wire			w_bus_valid;
	wire			w_bus_ready;
	wire	[7:0]	w_bus_wdata;
	wire	[7:0]	w_bus_rdata;
	wire			w_bus_rdata_en;

	wire			w_bus_vdp_ioreq;
	wire			w_bus_vdp_ready;
	wire	[7:0]	w_bus_vdp_rdata;
	wire			w_bus_vdp_rdata_en;

	wire			w_sdram_init_busy;

	// VDP <-> SDRAM VRAM bus
	wire	[22:2]	w_sdram_address;
	wire			w_sdram_write;
	wire			w_sdram_valid;
	wire			w_sdram_refresh;
	wire	[31:0]	w_sdram_wdata;
	wire	[3:0]	w_sdram_wdata_mask;
	wire	[31:0]	w_sdram_rdata;
	wire			w_sdram_rdata_en;

	// [MOD] Local wires for VDP VRAM bus (word address 17:0)
	wire	[17:0]	w_vram_address;
	wire	[31:0]	w_vram_wdata;
	wire	[31:0]	w_vram_rdata;
	wire			w_vram_valid;
	wire			w_vram_write;
	wire			w_vram_rdata_en;

	wire			w_video_de;
	wire			w_video_hs;
	wire			w_video_vs;
	wire	[7:0]	w_video_r;
	wire	[7:0]	w_video_g;
	wire	[7:0]	w_video_b;

	wire			w_pulse0;
	wire			w_pulse1;
	wire			w_pulse2;
	wire			w_pulse3;
	wire			w_pulse4;
	wire			w_pulse5;
	wire			w_pulse6;
	wire			w_pulse7;
	wire			w_wr;
	wire			w_sending;
	wire	[7:0]	w_red;
	wire	[7:0]	w_green;
	wire	[7:0]	w_blue;
	wire			w_int_n;

	assign slot_wait		= w_sdram_init_busy;
	assign oe_n				= 1'b0;

	always @( posedge clk85m ) begin
		ff_reset_n0		<= slot_reset_n;
		ff_reset_n1		<= ff_reset_n0;
		ff_reset_n2_1	<= ff_reset_n1;
		ff_reset_n2_2	<= ff_reset_n1;
	end

	assign reset_n	= ff_reset_n2_1;
	assign reset_n2	= ff_reset_n2_2;

	// --------------------------------------------------------------------
	//	clock
	// --------------------------------------------------------------------
	Gowin_rPLL u_pll (
		.clkout			( clk215m			),		//	output clkout	214.7727MHz
		.lock			( pll_lock215		),
		.clkin			( clk14m			)		//	input clkin		14.31818MHz
	);

	Gowin_rPLL2 u_pll2 (
		.clkout			( clk85m			),		//	output clkout	85.90908MHz
		.lock			( pll_lock85		),
		.clkoutp		( clk85m_n			),		//	output clkoutp	85.90908MHz (180deg phase shift)
		.clkin			( clk14m			)		//	input clkin		14.31818MHz
    );

	Gowin_CLKDIV u_clkdiv (
		.clkout			( clk42m			),		//	output clkout	42.95454MHz
		.hclkin			( clk85m			),		//	input hclkin	85.90908MHz
		.resetn			( pll_lock85		)		//	input resetn
	);

	// --------------------------------------------------------------------
	//	FullColor Intelligent LED
	// --------------------------------------------------------------------
	msx_slot u_msx_slot (
		.clk				( clk85m					),
		.initial_busy		( w_sdram_init_busy			),
		.p_slot_reset_n		( reset_n					),
		.p_slot_ioreq_n		( slot_iorq_n				),
		.p_slot_wr_n		( slot_wr_n					),
		.p_slot_rd_n		( slot_rd_n					),
		.p_slot_address		( slot_a					),
		.p_slot_data		( slot_d					),
		.p_slot_int			( slot_intr					),
		.p_slot_data_dir	( slot_data_dir				),
		.int_n				( w_int_n					),
		.bus_address		( w_bus_address				),
		.bus_ioreq			( w_bus_ioreq				),
		.bus_write			( w_bus_write				),
		.bus_valid			( w_bus_valid				),
		.bus_ready			( w_bus_ready				),
		.bus_wdata			( w_bus_wdata				),
		.bus_rdata			( w_bus_rdata				),
		.bus_rdata_en		( w_bus_rdata_en			),
		.dipsw				( dipsw[0]					)
	);

	assign w_bus_rdata		= ( w_bus_vdp_rdata_en		) ? w_bus_vdp_rdata: 8'hFF;
	assign w_bus_rdata_en	= w_bus_vdp_rdata_en;
	assign w_bus_ready		= w_bus_vdp_ready;

	// --------------------------------------------------------------------
	//	V9958 clone
	// --------------------------------------------------------------------
	vdp u_v9958 (
		.reset_n			( reset_n					),
		.clk				( clk85m					),
		.initial_busy		( w_sdram_init_busy			),
		.bus_address		( w_bus_address				),
		.bus_ioreq			( w_bus_ioreq				),
		.bus_write			( w_bus_write				),
		.bus_valid			( w_bus_valid				),
		.bus_ready			( w_bus_vdp_ready			),
		.bus_wdata			( w_bus_wdata				),
		.bus_rdata			( w_bus_vdp_rdata			),
		.bus_rdata_en		( w_bus_vdp_rdata_en		),
		.int_n				( w_int_n					),

		// [MOD] connect VDP VRAM bus to local wires
		.vram_address		( w_vram_address			),	// WORD address [17:0]
		.vram_write			( w_vram_write				),
		.vram_valid			( w_vram_valid				),
		.vram_wdata			( w_vram_wdata				),
		.vram_wdata_mask	( w_sdram_wdata_mask		),	// mask shared with SDRAM model
		.vram_rdata			( w_vram_rdata				),
		.vram_rdata_en		( w_vram_rdata_en			),
		.vram_refresh		( w_sdram_refresh			),

		.display_hs			( w_video_hs				),
		.display_vs			( w_video_vs				),
		.display_en			( w_video_de				),
		.display_r			( w_video_r					),
		.display_g			( w_video_g					),
		.display_b			( w_video_b					),
		.force_highspeed	( dipsw[1]					),
		.button				( button					),
		.pulse0				( w_pulse0					),
		.pulse1				( w_pulse1					),
		.pulse2				( w_pulse2					),
		.pulse3				( w_pulse3					),
		.pulse4				( w_pulse4					),
		.pulse5				( w_pulse5					),
		.pulse6				( w_pulse6					),
		.pulse7				( w_pulse7					)
	);

	// --------------------------------------------------------------------
	//	VRAM bus mapping
	// --------------------------------------------------------------------
	// Map VDP VRAM bus to SDRAM bus (original hardware behavior)
	// SDRAM address is 22:2, VDP provides 17:0 word address. Upper bits fixed to 0.
	assign w_sdram_address[22:18]	= 5'd0;
	assign w_sdram_address[17:2]	= w_vram_address;

	assign w_sdram_wdata			= w_vram_wdata;
	assign w_sdram_valid			= w_vram_valid;
	assign w_sdram_write			= w_vram_write;
// NOTE: do NOT create a circular assign between w_sdram_rdata_en and w_vram_rdata_en.
// The SDRAM model drives w_sdram_rdata_en; we expose that to the VDP by assigning
// w_vram_rdata_en := w_sdram_rdata_en (or to dbg_vram_rdata_en when requested).

// Use dbg_vram_* only when explicitly requested during Verilator runs.
// Default uses the SDRAM model (w_sdram_rdata).
`ifdef VERILATOR_DBGVRAM
  assign w_vram_rdata = dbg_vram_rdata;
  assign w_vram_rdata_en = dbg_vram_rdata_en;
`else
  assign w_vram_rdata = w_sdram_rdata;
  assign w_vram_rdata_en = w_sdram_rdata_en;
`endif


	// --------------------------------------------------------------------
	//	HDMI
	// --------------------------------------------------------------------
	DVI_TX_Top u_dvi (
		.I_rst_n			( reset_n2					),		//input I_rst_n
		.I_serial_clk		( clk215m					),		//input I_serial_clk
		.I_rgb_clk			( clk42m					),		//input I_rgb_clk
		.I_rgb_vs			( w_video_vs				),		//input I_rgb_vs
		.I_rgb_hs			( w_video_hs				),		//input I_rgb_hs
		.I_rgb_de			( w_video_de				),		//input I_rgb_de
		.I_rgb_r			( w_video_r					),		//input [7:0] I_rgb_r
		.I_rgb_g			( w_video_g					),		//input [7:0] I_rgb_g
		.I_rgb_b			( w_video_b					),		//input [7:0] I_rgb_b
		.O_tmds_clk_p		( tmds_clk_p				),		//output O_tmds_clk_p
		.O_tmds_clk_n		( tmds_clk_n				),		//output O_tmds_clk_n
		.O_tmds_data_p		( tmds_d_p					),		//output [2:0] O_tmds_data_p
		.O_tmds_data_n		( tmds_d_n					)		//output [2:0] O_tmds_data_n
	);

	// --------------------------------------------------------------------
	//	SDRAM
	// --------------------------------------------------------------------
	ip_sdram #(
		.FREQ				( 85_909_080				)		//	Hz
	) u_sdram (
		.reset_n			( reset_n					),
		.clk				( clk85m					),		//	85.90908MHz
		.clk_sdram			( clk85m_n					),
		.sdram_init_busy	( w_sdram_init_busy			),

		// [MOD] Use w_sdram_* signals that are already driven from VDP VRAM bus
		.bus_address		( w_sdram_address			),
		.bus_valid			( w_sdram_valid				),
		.bus_write			( w_sdram_write				),
		.bus_refresh		( w_sdram_refresh			),
		.bus_wdata			( w_sdram_wdata				),
		.bus_wdata_mask		( w_sdram_wdata_mask		),
		.bus_rdata			( w_sdram_rdata				),
		.bus_rdata_en		( w_sdram_rdata_en			),

		.O_sdram_clk		( O_sdram_clk				),
		.O_sdram_cke		( O_sdram_cke				),
		.O_sdram_cs_n		( O_sdram_cs_n				),		// chip select
		.O_sdram_ras_n		( O_sdram_ras_n				),		// row address select
		.O_sdram_cas_n		( O_sdram_cas_n				),		// columns address select
		.O_sdram_wen_n		( O_sdram_wen_n				),		// write enable
		.IO_sdram_dq		( IO_sdram_dq				),		// 32 bit bidirectional data bus
		.O_sdram_addr		( O_sdram_addr				),		// 11 bit multiplexed address bus
		.O_sdram_ba			( O_sdram_ba				),		// two banks
		.O_sdram_dqm		( O_sdram_dqm				)		// data mask
	);

	// --------------------------------------------------------------------
	//	Debug LED / Debugger (unchanged)
	// --------------------------------------------------------------------
	ip_ws2812_led u_led (
		.reset_n			( reset_n					),
		.clk				( clk85m					),
		.wr					( w_wr						),
		.sending			( w_sending					),
		.red				( w_red						),
		.green				( w_green					),
		.blue				( w_blue					),
		.ws2812_led			( ws2812_led				)
	);

	ip_debugger u_debugger (
		.reset_n			( reset_n					),
		.clk				( clk85m					),
		.pulse0				( w_pulse0					),
		.pulse1				( w_pulse1					),
		.pulse2				( w_pulse2					),
		.pulse3				( w_pulse3					),
		.pulse4				( w_pulse4					),
		.pulse5				( w_pulse5					),
		.pulse6				( w_pulse6					),
		.pulse7				( w_pulse7					),
		.wr					( w_wr						),
		.sending			( w_sending					),
		.red				( w_red						),
		.green				( w_green					),
		.blue				( w_blue					)
	);

	// --------------------------------------------------------------------
	// [MOD] Export VRAM bus for Verilator/C++ wrapper
	// --------------------------------------------------------------------
	assign dbg_vram_address	= w_vram_address;
	assign dbg_vram_wdata	= w_vram_wdata;
	assign dbg_vram_valid	= w_vram_valid;
	assign dbg_vram_write	= w_vram_write;
	assign dbg_vram_rdata_en= w_vram_rdata_en;

	// --------------------------------------------------------------------
	// [MOD] Export VIDEO Out for Verilator/C++ wrapper
	// --------------------------------------------------------------------
    assign display_hs = w_video_hs;
    assign display_vs = w_video_vs;
    assign display_en = w_video_de;
    assign display_r  = w_video_r;
    assign display_g  = w_video_g;
    assign display_b  = w_video_b;
	
// --------------------------------------------------------------------
// Debug monitors (Verilator only)
//
// These prints help confirm the rdata_en path:
//  - SDRAM model asserts w_sdram_rdata_en
//  - top should observe w_sdram_rdata_en
//  - vdp_vram_interface should see vram_rdata_en (which is driven from w_sdram_rdata_en)
// Guarded by `ifdef VERILATOR to avoid synthesis impacts.
// --------------------------------------------------------------------
`ifdef VERILATOR
	reg prev_sdram_rdata_en;
	reg prev_vram_rdata_en;
	always @(posedge clk85m) begin
		if (!reset_n) begin
			prev_sdram_rdata_en <= 1'b0;
			prev_vram_rdata_en  <= 1'b0;
		end else begin
			prev_sdram_rdata_en <= w_sdram_rdata_en;
			prev_vram_rdata_en  <= w_vram_rdata_en;
		end
	end
`endif

endmodule